module RegisterFile(regA, regB, Destreg, Data, en, contRegA, contRegB);
  input [2:0] regA, regB, Destreg;
  input en;
  input [31:0] Data;
  output [31:0] contRegA, contRegB;

  
endmodule