module Decoder()

endmodule