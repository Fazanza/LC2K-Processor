module Adder(in1, in2, outVal);
  input [7:0] in1, in2;
  output [15:0] outVal;

  assign outVal = in1, in2;
endmodule