module Processor(clk);
  input clk;

  reg a;
  always @(posedge clk) begin
    
  end
endmodule