module Processor(clk);
  input clk;

  always @(posedge clk) begin
    
  end
endmodule